module top(
    input wire [7:9] i_select, hello_there_haha
    input i_clk0,
    input i_clk1,
    output o_clk
    );



endmodule
